module Instruction_Memory #(parameter ADDRESS_WIDTH = 20, parameter DATA_WIDTH = 32)
(
    input Enable,
    input [ADDRESS_WIDTH - 1 : 0] Address,

    output [DATA_WIDTH - 1 : 0] Data
);

    reg [DATA_WIDTH - 1 : 0] Memory [$pow(2, ADDRESS_WIDTH) - 1 : 0];

    initial
    begin
		Memory[0]	=	32'h4e583111;
		Memory[1]	=	32'h49c30922;
		Memory[2]	=	32'h42beee82;
		Memory[3]	=	32'he9406ab1;
		Memory[4]	=	32'h80a545c5;
		Memory[5]	=	32'h9bd8d943;
		Memory[6]	=	32'h99f4ffb7;
		Memory[7]	=	32'hf325f246;
		Memory[8]	=	32'h6e8da1ce;
		Memory[9]	=	32'h1be20f9f;
		Memory[10]	=	32'h992c5e1b;
		Memory[11]	=	32'h419f421b;
		Memory[12]	=	32'h64c0bfba;
		Memory[13]	=	32'h8234b878;
		Memory[14]	=	32'h49aa8b3f;
		Memory[15]	=	32'h82d865c1;
		Memory[16]	=	32'hce61e8c1;
		Memory[17]	=	32'h93594ba0;
		Memory[18]	=	32'h508f936;
		Memory[19]	=	32'hb088ced6;
		Memory[20]	=	32'hb2ba6cd5;
		Memory[21]	=	32'h6b069ff;
		Memory[22]	=	32'hf23f005f;
		Memory[23]	=	32'h9adec517;
		Memory[24]	=	32'hfdaf238;
		Memory[25]	=	32'h64d4dcb2;
		Memory[26]	=	32'hb6790da2;
		Memory[27]	=	32'hbe423970;
		Memory[28]	=	32'h415ac756;
		Memory[29]	=	32'hbb79e6ed;
		Memory[30]	=	32'hd2c08fe2;
		Memory[31]	=	32'h3eec7c09;
		Memory[32]	=	32'h6033af0;
		Memory[33]	=	32'h529583a6;
		Memory[34]	=	32'h27c28045;
		Memory[35]	=	32'hf6862995;
		Memory[36]	=	32'h29e39259;
		Memory[37]	=	32'h3e8fe397;
		Memory[38]	=	32'h745c53d3;
		Memory[39]	=	32'h5b319790;
		Memory[40]	=	32'h5811ceb8;
		Memory[41]	=	32'hd51c9c3;
		Memory[42]	=	32'h25d3905c;
		Memory[43]	=	32'h4576208d;
		Memory[44]	=	32'h8e22de38;
		Memory[45]	=	32'he3d75f02;
		Memory[46]	=	32'h5cc6bbef;
		Memory[47]	=	32'ha4311f45;
		Memory[48]	=	32'h18984958;
		Memory[49]	=	32'h58afe0c;
		Memory[50]	=	32'h61d6f5e8;
		Memory[51]	=	32'h9ff9c796;
		Memory[52]	=	32'h698e5431;
		Memory[53]	=	32'hc3c726e;
		Memory[54]	=	32'h7ec48a8e;
		Memory[55]	=	32'h51f8ca32;
		Memory[56]	=	32'hff5cc0d4;
		Memory[57]	=	32'hee76dfeb;
		Memory[58]	=	32'hbf1b8463;
		Memory[59]	=	32'h3054651e;
		Memory[60]	=	32'h73f961c9;
		Memory[61]	=	32'h26b19349;
		Memory[62]	=	32'hba1b5043;
		Memory[63]	=	32'hbe18d8db;
		Memory[64]	=	32'h213f2395;
		Memory[65]	=	32'h7a8b5336;
		Memory[66]	=	32'hb552f1a;
		Memory[67]	=	32'h746c335b;
		Memory[68]	=	32'h9a86a55a;
		Memory[69]	=	32'h1cb50242;
		Memory[70]	=	32'hef54aae8;
		Memory[71]	=	32'heaffdea0;
		Memory[72]	=	32'h17f1327e;
		Memory[73]	=	32'hcce54048;
		Memory[74]	=	32'h8b023acb;
		Memory[75]	=	32'hbd99d40c;
		Memory[76]	=	32'ha4621ee0;
		Memory[77]	=	32'hd522cb08;
		Memory[78]	=	32'h409a283c;
		Memory[79]	=	32'h8cf11655;
		Memory[80]	=	32'h83440f4e;
		Memory[81]	=	32'he0737a40;
		Memory[82]	=	32'he4aaf8bb;
		Memory[83]	=	32'hc0fef5e6;
		Memory[84]	=	32'h45ce770;
		Memory[85]	=	32'he45410f5;
		Memory[86]	=	32'h1bb569d9;
		Memory[87]	=	32'h8d771f;
		Memory[88]	=	32'hf49870cd;
		Memory[89]	=	32'h6365464e;
		Memory[90]	=	32'hf3f72df8;
		Memory[91]	=	32'h375bd03d;
		Memory[92]	=	32'h43d70239;
		Memory[93]	=	32'h62f03d6a;
		Memory[94]	=	32'hbbb1019f;
		Memory[95]	=	32'h9bab63a1;
		Memory[96]	=	32'h7138f258;
		Memory[97]	=	32'ha0a621b0;
		Memory[98]	=	32'hb7043507;
		Memory[99]	=	32'hc118244c;
    end

    assign Data = Enable ? Memory[Address] : 'bz;
endmodule
